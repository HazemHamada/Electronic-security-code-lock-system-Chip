LIBRARY sxlib_ModelSim;

entity sdetj_b_l is
   port (
      vdd     : in      bit;
      clk     : in      bit;
      vss     : in      bit;
      reset   : in      bit;
      daytime : in      bit;
      code    : in      bit_vector(3 downto 0);
      door    : out     bit;
      alarm   : out     bit
 );
end sdetj_b_l;

architecture structural of sdetj_b_l is
Component a4_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      i3  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component an12_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component inv_x2
   port (
      i   : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component no4_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      i3  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component oa22_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component xr2_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component ao22_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component no2_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component a2_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component o4_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      i3  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component nao22_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component o3_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component on12_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component o2_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component na3_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component sff1_x4
   port (
      ck  : in      bit;
      i   : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component no3_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component na4_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      i3  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component na2_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

signal dacs_cs        : bit_vector( 2 downto 0);
signal not_code       : bit_vector( 3 downto 1);
signal not_dacs_cs    : bit_vector( 2 downto 1);
signal xr2_x1_sig     : bit;
signal on12_x1_sig    : bit;
signal oa22_x2_sig    : bit;
signal o4_x2_sig      : bit;
signal o3_x2_sig      : bit;
signal o3_x2_3_sig    : bit;
signal o3_x2_2_sig    : bit;
signal o2_x2_sig      : bit;
signal not_reset      : bit;
signal not_aux9       : bit;
signal not_aux8       : bit;
signal not_aux15      : bit;
signal not_aux13      : bit;
signal not_aux12      : bit;
signal not_aux11      : bit;
signal not_aux1       : bit;
signal not_aux0       : bit;
signal no2_x1_sig     : bit;
signal nao22_x1_sig   : bit;
signal nao22_x1_2_sig : bit;
signal na4_x1_sig     : bit;
signal na3_x1_sig     : bit;
signal na3_x1_5_sig   : bit;
signal na3_x1_4_sig   : bit;
signal na3_x1_3_sig   : bit;
signal na3_x1_2_sig   : bit;
signal na2_x1_sig     : bit;
signal na2_x1_3_sig   : bit;
signal na2_x1_2_sig   : bit;
signal inv_x2_sig     : bit;
signal aux4           : bit;
signal ao22_x2_sig    : bit;
signal a4_x2_sig      : bit;
signal a2_x2_sig      : bit;

begin

not_aux11_ins : o2_x2
   port map (
      i0  => reset,
      i1  => dacs_cs(2),
      q   => not_aux11,
      vdd => vdd,
      vss => vss
   );

na2_x1_ins : na2_x1
   port map (
      i0  => not_aux12,
      i1  => dacs_cs(1),
      nq  => na2_x1_sig,
      vdd => vdd,
      vss => vss
   );

na2_x1_2_ins : na2_x1
   port map (
      i0  => not_aux9,
      i1  => dacs_cs(1),
      nq  => na2_x1_2_sig,
      vdd => vdd,
      vss => vss
   );

not_aux15_ins : na3_x1
   port map (
      i0  => na2_x1_2_sig,
      i1  => dacs_cs(0),
      i2  => na2_x1_sig,
      nq  => not_aux15,
      vdd => vdd,
      vss => vss
   );

not_aux0_ins : o2_x2
   port map (
      i0  => dacs_cs(0),
      i1  => dacs_cs(1),
      q   => not_aux0,
      vdd => vdd,
      vss => vss
   );

a4_x2_ins : a4_x2
   port map (
      i0  => not_reset,
      i1  => daytime,
      i2  => code(2),
      i3  => code(3),
      q   => a4_x2_sig,
      vdd => vdd,
      vss => vss
   );

not_aux8_ins : on12_x1
   port map (
      i0  => a4_x2_sig,
      i1  => not_aux1,
      q   => not_aux8,
      vdd => vdd,
      vss => vss
   );

not_aux12_ins : o2_x2
   port map (
      i0  => code(3),
      i1  => not_code(2),
      q   => not_aux12,
      vdd => vdd,
      vss => vss
   );

not_dacs_cs_2_ins : inv_x2
   port map (
      i   => dacs_cs(2),
      nq  => not_dacs_cs(2),
      vdd => vdd,
      vss => vss
   );

not_aux9_ins : o2_x2
   port map (
      i0  => code(0),
      i1  => not_code(1),
      q   => not_aux9,
      vdd => vdd,
      vss => vss
   );

not_dacs_cs_1_ins : inv_x2
   port map (
      i   => dacs_cs(1),
      nq  => not_dacs_cs(1),
      vdd => vdd,
      vss => vss
   );

not_aux13_ins : an12_x1
   port map (
      i0  => aux4,
      i1  => not_reset,
      q   => not_aux13,
      vdd => vdd,
      vss => vss
   );

not_aux1_ins : on12_x1
   port map (
      i0  => code(0),
      i1  => code(1),
      q   => not_aux1,
      vdd => vdd,
      vss => vss
   );

not_reset_ins : inv_x2
   port map (
      i   => reset,
      nq  => not_reset,
      vdd => vdd,
      vss => vss
   );

not_code_3_ins : inv_x2
   port map (
      i   => code(3),
      nq  => not_code(3),
      vdd => vdd,
      vss => vss
   );

not_code_2_ins : inv_x2
   port map (
      i   => code(2),
      nq  => not_code(2),
      vdd => vdd,
      vss => vss
   );

not_code_1_ins : inv_x2
   port map (
      i   => code(1),
      nq  => not_code(1),
      vdd => vdd,
      vss => vss
   );

inv_x2_ins : inv_x2
   port map (
      i   => daytime,
      nq  => inv_x2_sig,
      vdd => vdd,
      vss => vss
   );

aux4_ins : no4_x1
   port map (
      i0  => not_code(2),
      i1  => inv_x2_sig,
      i2  => not_aux1,
      i3  => not_code(3),
      nq  => aux4,
      vdd => vdd,
      vss => vss
   );

na2_x1_3_ins : na2_x1
   port map (
      i0  => dacs_cs(0),
      i1  => dacs_cs(2),
      nq  => na2_x1_3_sig,
      vdd => vdd,
      vss => vss
   );

o3_x2_ins : o3_x2
   port map (
      i0  => code(3),
      i1  => code(2),
      i2  => not_aux9,
      q   => o3_x2_sig,
      vdd => vdd,
      vss => vss
   );

oa22_x2_ins : oa22_x2
   port map (
      i0  => not_dacs_cs(1),
      i1  => o3_x2_sig,
      i2  => na2_x1_3_sig,
      q   => oa22_x2_sig,
      vdd => vdd,
      vss => vss
   );

xr2_x1_ins : xr2_x1
   port map (
      i0  => dacs_cs(1),
      i1  => dacs_cs(0),
      q   => xr2_x1_sig,
      vdd => vdd,
      vss => vss
   );

nao22_x1_ins : nao22_x1
   port map (
      i0  => not_aux1,
      i1  => not_aux12,
      i2  => dacs_cs(1),
      nq  => nao22_x1_sig,
      vdd => vdd,
      vss => vss
   );

na3_x1_2_ins : na3_x1
   port map (
      i0  => not_dacs_cs(2),
      i1  => nao22_x1_sig,
      i2  => xr2_x1_sig,
      nq  => na3_x1_2_sig,
      vdd => vdd,
      vss => vss
   );

na3_x1_ins : na3_x1
   port map (
      i0  => not_aux13,
      i1  => na3_x1_2_sig,
      i2  => oa22_x2_sig,
      nq  => na3_x1_sig,
      vdd => vdd,
      vss => vss
   );

dacs_cs_0_ins : sff1_x4
   port map (
      ck  => clk,
      i   => na3_x1_sig,
      q   => dacs_cs(0),
      vdd => vdd,
      vss => vss
   );

ao22_x2_ins : ao22_x2
   port map (
      i0  => not_aux15,
      i1  => not_aux11,
      i2  => not_aux8,
      q   => ao22_x2_sig,
      vdd => vdd,
      vss => vss
   );

o3_x2_2_ins : o3_x2
   port map (
      i0  => code(0),
      i1  => code(1),
      i2  => not_aux0,
      q   => o3_x2_2_sig,
      vdd => vdd,
      vss => vss
   );

no2_x1_ins : no2_x1
   port map (
      i0  => code(0),
      i1  => not_code(1),
      nq  => no2_x1_sig,
      vdd => vdd,
      vss => vss
   );

na3_x1_3_ins : na3_x1
   port map (
      i0  => no2_x1_sig,
      i1  => dacs_cs(0),
      i2  => not_dacs_cs(1),
      nq  => na3_x1_3_sig,
      vdd => vdd,
      vss => vss
   );

a2_x2_ins : a2_x2
   port map (
      i0  => na3_x1_3_sig,
      i1  => o3_x2_2_sig,
      q   => a2_x2_sig,
      vdd => vdd,
      vss => vss
   );

o4_x2_ins : o4_x2
   port map (
      i0  => reset,
      i1  => code(3),
      i2  => code(2),
      i3  => not_dacs_cs(2),
      q   => o4_x2_sig,
      vdd => vdd,
      vss => vss
   );

nao22_x1_2_ins : nao22_x1
   port map (
      i0  => o4_x2_sig,
      i1  => a2_x2_sig,
      i2  => ao22_x2_sig,
      nq  => nao22_x1_2_sig,
      vdd => vdd,
      vss => vss
   );

dacs_cs_1_ins : sff1_x4
   port map (
      ck  => clk,
      i   => nao22_x1_2_sig,
      q   => dacs_cs(1),
      vdd => vdd,
      vss => vss
   );

o3_x2_3_ins : o3_x2
   port map (
      i0  => not_code(3),
      i1  => code(2),
      i2  => not_aux9,
      q   => o3_x2_3_sig,
      vdd => vdd,
      vss => vss
   );

on12_x1_ins : on12_x1
   port map (
      i0  => o3_x2_3_sig,
      i1  => dacs_cs(0),
      q   => on12_x1_sig,
      vdd => vdd,
      vss => vss
   );

na3_x1_5_ins : na3_x1
   port map (
      i0  => dacs_cs(2),
      i1  => dacs_cs(1),
      i2  => on12_x1_sig,
      nq  => na3_x1_5_sig,
      vdd => vdd,
      vss => vss
   );

o2_x2_ins : o2_x2
   port map (
      i0  => not_aux15,
      i1  => dacs_cs(2),
      q   => o2_x2_sig,
      vdd => vdd,
      vss => vss
   );

na3_x1_4_ins : na3_x1
   port map (
      i0  => not_aux13,
      i1  => o2_x2_sig,
      i2  => na3_x1_5_sig,
      nq  => na3_x1_4_sig,
      vdd => vdd,
      vss => vss
   );

dacs_cs_2_ins : sff1_x4
   port map (
      ck  => clk,
      i   => na3_x1_4_sig,
      q   => dacs_cs(2),
      vdd => vdd,
      vss => vss
   );

alarm_ins : no3_x1
   port map (
      i0  => aux4,
      i1  => not_aux11,
      i2  => not_aux0,
      nq  => alarm,
      vdd => vdd,
      vss => vss
   );

na4_x1_ins : na4_x1
   port map (
      i0  => dacs_cs(2),
      i1  => not_reset,
      i2  => dacs_cs(0),
      i3  => dacs_cs(1),
      nq  => na4_x1_sig,
      vdd => vdd,
      vss => vss
   );

door_ins : na2_x1
   port map (
      i0  => not_aux8,
      i1  => na4_x1_sig,
      nq  => door,
      vdd => vdd,
      vss => vss
   );


end structural;
